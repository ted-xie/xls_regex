module __donut__donut(
  input wire clk,
  input wire [127:0] stream,
  output wire [15:0] out
);
  function automatic [0:0] bit_slice_update_w1_1b_1b (input reg [0:0] to_update, input reg [0:0] start, input reg [0:0] update_value);
    begin
      bit_slice_update_w1_1b_1b = start >= 1'h1 ? to_update : update_value << start | ~(1'h1 << start) & to_update;
    end
  endfunction
  wire [255:0] literal_59710;
  assign literal_59710 = {1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h1, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0};
  wire [7:0] stream_unflattened[16];
  assign stream_unflattened[0] = stream[127:120];
  assign stream_unflattened[1] = stream[119:112];
  assign stream_unflattened[2] = stream[111:104];
  assign stream_unflattened[3] = stream[103:96];
  assign stream_unflattened[4] = stream[95:88];
  assign stream_unflattened[5] = stream[87:80];
  assign stream_unflattened[6] = stream[79:72];
  assign stream_unflattened[7] = stream[71:64];
  assign stream_unflattened[8] = stream[63:56];
  assign stream_unflattened[9] = stream[55:48];
  assign stream_unflattened[10] = stream[47:40];
  assign stream_unflattened[11] = stream[39:32];
  assign stream_unflattened[12] = stream[31:24];
  assign stream_unflattened[13] = stream[23:16];
  assign stream_unflattened[14] = stream[15:8];
  assign stream_unflattened[15] = stream[7:0];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_stream[15:0];
  always_ff @ (posedge clk) begin
    //p0_stream <= stream_unflattened;
    p0_stream[0] <= stream_unflattened[0];
    p0_stream[1] <= stream_unflattened[1];
    p0_stream[2] <= stream_unflattened[2];
    p0_stream[3] <= stream_unflattened[3];
    p0_stream[4] <= stream_unflattened[4];
    p0_stream[5] <= stream_unflattened[5];
    p0_stream[6] <= stream_unflattened[6];
    p0_stream[7] <= stream_unflattened[7];
    p0_stream[8] <= stream_unflattened[8];
    p0_stream[9] <= stream_unflattened[9];
    p0_stream[10] <= stream_unflattened[10];
    p0_stream[11] <= stream_unflattened[11];
    p0_stream[12] <= stream_unflattened[12];
    p0_stream[13] <= stream_unflattened[13];
    p0_stream[14] <= stream_unflattened[14];
    p0_stream[15] <= stream_unflattened[15];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_ch_comb;
  wire [7:0] p1_ch__1_comb;
  wire [7:0] p1_ch__2_comb;
  wire [7:0] p1_ch__3_comb;
  wire [7:0] p1_ch__4_comb;
  wire [7:0] p1_ch__5_comb;
  wire [7:0] p1_ch__6_comb;
  wire [7:0] p1_ch__7_comb;
  wire [7:0] p1_ch__8_comb;
  wire [7:0] p1_ch__9_comb;
  wire [7:0] p1_ch__10_comb;
  wire [7:0] p1_ch__11_comb;
  wire [7:0] p1_ch__12_comb;
  wire [7:0] p1_ch__13_comb;
  wire [7:0] p1_ch__14_comb;
  wire [7:0] p1_ch__15_comb;
  wire p1_result_i__4_comb;
  wire p1_result_i__145_comb;
  wire p1_accept_ch__10_comb;
  wire p1_result_i__149_comb;
  wire p1_result_i__150_comb;
  wire p1_accept_ch__29_comb;
  wire p1_result_i__154_comb;
  wire p1_result_i__155_comb;
  wire p1_accept_ch__45_comb;
  wire p1_result_i__159_comb;
  wire p1_result_i__160_comb;
  wire p1_accept_ch__61_comb;
  wire p1_result_i__164_comb;
  wire p1_result_i__165_comb;
  wire p1_accept_ch__77_comb;
  wire p1_result_i__169_comb;
  wire p1_result_i__170_comb;
  wire p1_accept_ch__93_comb;
  wire p1_result_i__174_comb;
  wire p1_result_i__175_comb;
  wire p1_accept_ch__109_comb;
  wire p1_result_i__179_comb;
  wire p1_result_i__180_comb;
  wire p1_accept_ch__125_comb;
  wire p1_result_i__184_comb;
  wire p1_result_i__185_comb;
  wire p1_accept_ch__141_comb;
  wire p1_result_i__189_comb;
  wire p1_result_i__190_comb;
  wire p1_accept_ch__157_comb;
  wire p1_result_i__194_comb;
  wire p1_result_i__195_comb;
  wire p1_accept_ch__173_comb;
  wire p1_result_i__199_comb;
  wire p1_result_i__200_comb;
  wire p1_accept_ch__189_comb;
  wire p1_result_i__204_comb;
  wire p1_result_i__205_comb;
  wire p1_accept_ch__205_comb;
  wire p1_result_i__209_comb;
  wire p1_result_i__210_comb;
  wire p1_accept_ch__221_comb;
  wire p1_result_i__214_comb;
  wire p1_result_i__215_comb;
  wire p1_accept_ch__237_comb;
  wire p1_result_i__219_comb;
  wire p1_result_i__220_comb;
  wire p1_accept_ch__253_comb;
  wire p1_result_i__146_comb;
  wire p1_result_i__5_comb;
  wire p1_result_i__151_comb;
  wire p1_result_i__14_comb;
  wire p1_result_i__156_comb;
  wire p1_result_i__23_comb;
  wire p1_result_i__161_comb;
  wire p1_result_i__32_comb;
  wire p1_result_i__166_comb;
  wire p1_result_i__41_comb;
  wire p1_result_i__171_comb;
  wire p1_result_i__50_comb;
  wire p1_result_i__176_comb;
  wire p1_result_i__59_comb;
  wire p1_result_i__181_comb;
  wire p1_result_i__68_comb;
  wire p1_result_i__186_comb;
  wire p1_result_i__77_comb;
  wire p1_result_i__191_comb;
  wire p1_result_i__86_comb;
  wire p1_result_i__196_comb;
  wire p1_result_i__95_comb;
  wire p1_result_i__201_comb;
  wire p1_result_i__104_comb;
  wire p1_result_i__206_comb;
  wire p1_result_i__113_comb;
  wire p1_result_i__211_comb;
  wire p1_result_i__122_comb;
  wire p1_result_i__216_comb;
  wire p1_result_i__131_comb;
  wire p1_result_i__221_comb;
  wire p1_result_i__140_comb;
  wire p1_result_i__147_comb;
  wire p1_result_i__6_comb;
  wire p1_result_i__152_comb;
  wire p1_result_i__15_comb;
  wire p1_result_i__157_comb;
  wire p1_result_i__24_comb;
  wire p1_result_i__162_comb;
  wire p1_result_i__33_comb;
  wire p1_result_i__167_comb;
  wire p1_result_i__42_comb;
  wire p1_result_i__172_comb;
  wire p1_result_i__51_comb;
  wire p1_result_i__177_comb;
  wire p1_result_i__60_comb;
  wire p1_result_i__182_comb;
  wire p1_result_i__69_comb;
  wire p1_result_i__187_comb;
  wire p1_result_i__78_comb;
  wire p1_result_i__192_comb;
  wire p1_result_i__87_comb;
  wire p1_result_i__197_comb;
  wire p1_result_i__96_comb;
  wire p1_result_i__202_comb;
  wire p1_result_i__105_comb;
  wire p1_result_i__207_comb;
  wire p1_result_i__114_comb;
  wire p1_result_i__212_comb;
  wire p1_result_i__123_comb;
  wire p1_result_i__217_comb;
  wire p1_result_i__132_comb;
  wire p1_result_i__222_comb;
  wire p1_result_i__141_comb;
  wire p1_result_i__148_comb;
  wire p1_result_i__7_comb;
  wire p1_result_i__153_comb;
  wire p1_result_i__16_comb;
  wire p1_result_i__158_comb;
  wire p1_result_i__25_comb;
  wire p1_result_i__163_comb;
  wire p1_result_i__34_comb;
  wire p1_result_i__168_comb;
  wire p1_result_i__43_comb;
  wire p1_result_i__173_comb;
  wire p1_result_i__52_comb;
  wire p1_result_i__178_comb;
  wire p1_result_i__61_comb;
  wire p1_result_i__183_comb;
  wire p1_result_i__70_comb;
  wire p1_result_i__188_comb;
  wire p1_result_i__79_comb;
  wire p1_result_i__193_comb;
  wire p1_result_i__88_comb;
  wire p1_result_i__198_comb;
  wire p1_result_i__97_comb;
  wire p1_result_i__203_comb;
  wire p1_result_i__106_comb;
  wire p1_result_i__208_comb;
  wire p1_result_i__115_comb;
  wire p1_result_i__213_comb;
  wire p1_result_i__124_comb;
  wire p1_result_i__218_comb;
  wire p1_result_i__133_comb;
  wire p1_result_i__223_comb;
  wire p1_result_i__142_comb;
  wire p1_result_i__8_comb;
  wire p1_result_i__17_comb;
  wire p1_result_i__26_comb;
  wire p1_result_i__35_comb;
  wire p1_result_i__44_comb;
  wire p1_result_i__53_comb;
  wire p1_result_i__62_comb;
  wire p1_result_i__71_comb;
  wire p1_result_i__80_comb;
  wire p1_result_i__89_comb;
  wire p1_result_i__98_comb;
  wire p1_result_i__107_comb;
  wire p1_result_i__116_comb;
  wire p1_result_i__125_comb;
  wire p1_result_i__134_comb;
  wire p1_result_i__143_comb;
  wire [15:0] p1_result__16_comb;
  assign p1_ch_comb = p0_stream[32'h0000_0000];
  assign p1_ch__1_comb = p0_stream[32'h0000_0001];
  assign p1_ch__2_comb = p0_stream[32'h0000_0002];
  assign p1_ch__3_comb = p0_stream[32'h0000_0003];
  assign p1_ch__4_comb = p0_stream[32'h0000_0004];
  assign p1_ch__5_comb = p0_stream[32'h0000_0005];
  assign p1_ch__6_comb = p0_stream[32'h0000_0006];
  assign p1_ch__7_comb = p0_stream[32'h0000_0007];
  assign p1_ch__8_comb = p0_stream[32'h0000_0008];
  assign p1_ch__9_comb = p0_stream[32'h0000_0009];
  assign p1_ch__10_comb = p0_stream[32'h0000_000a];
  assign p1_ch__11_comb = p0_stream[32'h0000_000b];
  assign p1_ch__12_comb = p0_stream[32'h0000_000c];
  assign p1_ch__13_comb = p0_stream[32'h0000_000d];
  assign p1_ch__14_comb = p0_stream[32'h0000_000e];
  assign p1_ch__15_comb = p0_stream[32'h0000_000f];
  assign p1_result_i__4_comb = 1'h0;
  assign p1_result_i__145_comb = 1'h0;
  assign p1_accept_ch__10_comb = literal_59710[p1_ch_comb];
  assign p1_result_i__149_comb = 1'h0;
  assign p1_result_i__150_comb = 1'h0;
  assign p1_accept_ch__29_comb = literal_59710[p1_ch__1_comb];
  assign p1_result_i__154_comb = 1'h0;
  assign p1_result_i__155_comb = 1'h0;
  assign p1_accept_ch__45_comb = literal_59710[p1_ch__2_comb];
  assign p1_result_i__159_comb = 1'h0;
  assign p1_result_i__160_comb = 1'h0;
  assign p1_accept_ch__61_comb = literal_59710[p1_ch__3_comb];
  assign p1_result_i__164_comb = 1'h0;
  assign p1_result_i__165_comb = 1'h0;
  assign p1_accept_ch__77_comb = literal_59710[p1_ch__4_comb];
  assign p1_result_i__169_comb = 1'h0;
  assign p1_result_i__170_comb = 1'h0;
  assign p1_accept_ch__93_comb = literal_59710[p1_ch__5_comb];
  assign p1_result_i__174_comb = 1'h0;
  assign p1_result_i__175_comb = 1'h0;
  assign p1_accept_ch__109_comb = literal_59710[p1_ch__6_comb];
  assign p1_result_i__179_comb = 1'h0;
  assign p1_result_i__180_comb = 1'h0;
  assign p1_accept_ch__125_comb = literal_59710[p1_ch__7_comb];
  assign p1_result_i__184_comb = 1'h0;
  assign p1_result_i__185_comb = 1'h0;
  assign p1_accept_ch__141_comb = literal_59710[p1_ch__8_comb];
  assign p1_result_i__189_comb = 1'h0;
  assign p1_result_i__190_comb = 1'h0;
  assign p1_accept_ch__157_comb = literal_59710[p1_ch__9_comb];
  assign p1_result_i__194_comb = 1'h0;
  assign p1_result_i__195_comb = 1'h0;
  assign p1_accept_ch__173_comb = literal_59710[p1_ch__10_comb];
  assign p1_result_i__199_comb = 1'h0;
  assign p1_result_i__200_comb = 1'h0;
  assign p1_accept_ch__189_comb = literal_59710[p1_ch__11_comb];
  assign p1_result_i__204_comb = 1'h0;
  assign p1_result_i__205_comb = 1'h0;
  assign p1_accept_ch__205_comb = literal_59710[p1_ch__12_comb];
  assign p1_result_i__209_comb = 1'h0;
  assign p1_result_i__210_comb = 1'h0;
  assign p1_accept_ch__221_comb = literal_59710[p1_ch__13_comb];
  assign p1_result_i__214_comb = 1'h0;
  assign p1_result_i__215_comb = 1'h0;
  assign p1_accept_ch__237_comb = literal_59710[p1_ch__14_comb];
  assign p1_result_i__219_comb = 1'h0;
  assign p1_result_i__220_comb = 1'h0;
  assign p1_accept_ch__253_comb = literal_59710[p1_ch__15_comb];
  assign p1_result_i__146_comb = 1'h0;
  assign p1_result_i__5_comb = bit_slice_update_w1_1b_1b(p1_result_i__4_comb, p1_result_i__145_comb, p1_accept_ch__10_comb);
  assign p1_result_i__151_comb = 1'h0;
  assign p1_result_i__14_comb = bit_slice_update_w1_1b_1b(p1_result_i__149_comb, p1_result_i__150_comb, p1_accept_ch__29_comb);
  assign p1_result_i__156_comb = 1'h0;
  assign p1_result_i__23_comb = bit_slice_update_w1_1b_1b(p1_result_i__154_comb, p1_result_i__155_comb, p1_accept_ch__45_comb);
  assign p1_result_i__161_comb = 1'h0;
  assign p1_result_i__32_comb = bit_slice_update_w1_1b_1b(p1_result_i__159_comb, p1_result_i__160_comb, p1_accept_ch__61_comb);
  assign p1_result_i__166_comb = 1'h0;
  assign p1_result_i__41_comb = bit_slice_update_w1_1b_1b(p1_result_i__164_comb, p1_result_i__165_comb, p1_accept_ch__77_comb);
  assign p1_result_i__171_comb = 1'h0;
  assign p1_result_i__50_comb = bit_slice_update_w1_1b_1b(p1_result_i__169_comb, p1_result_i__170_comb, p1_accept_ch__93_comb);
  assign p1_result_i__176_comb = 1'h0;
  assign p1_result_i__59_comb = bit_slice_update_w1_1b_1b(p1_result_i__174_comb, p1_result_i__175_comb, p1_accept_ch__109_comb);
  assign p1_result_i__181_comb = 1'h0;
  assign p1_result_i__68_comb = bit_slice_update_w1_1b_1b(p1_result_i__179_comb, p1_result_i__180_comb, p1_accept_ch__125_comb);
  assign p1_result_i__186_comb = 1'h0;
  assign p1_result_i__77_comb = bit_slice_update_w1_1b_1b(p1_result_i__184_comb, p1_result_i__185_comb, p1_accept_ch__141_comb);
  assign p1_result_i__191_comb = 1'h0;
  assign p1_result_i__86_comb = bit_slice_update_w1_1b_1b(p1_result_i__189_comb, p1_result_i__190_comb, p1_accept_ch__157_comb);
  assign p1_result_i__196_comb = 1'h0;
  assign p1_result_i__95_comb = bit_slice_update_w1_1b_1b(p1_result_i__194_comb, p1_result_i__195_comb, p1_accept_ch__173_comb);
  assign p1_result_i__201_comb = 1'h0;
  assign p1_result_i__104_comb = bit_slice_update_w1_1b_1b(p1_result_i__199_comb, p1_result_i__200_comb, p1_accept_ch__189_comb);
  assign p1_result_i__206_comb = 1'h0;
  assign p1_result_i__113_comb = bit_slice_update_w1_1b_1b(p1_result_i__204_comb, p1_result_i__205_comb, p1_accept_ch__205_comb);
  assign p1_result_i__211_comb = 1'h0;
  assign p1_result_i__122_comb = bit_slice_update_w1_1b_1b(p1_result_i__209_comb, p1_result_i__210_comb, p1_accept_ch__221_comb);
  assign p1_result_i__216_comb = 1'h0;
  assign p1_result_i__131_comb = bit_slice_update_w1_1b_1b(p1_result_i__214_comb, p1_result_i__215_comb, p1_accept_ch__237_comb);
  assign p1_result_i__221_comb = 1'h0;
  assign p1_result_i__140_comb = bit_slice_update_w1_1b_1b(p1_result_i__219_comb, p1_result_i__220_comb, p1_accept_ch__253_comb);
  assign p1_result_i__147_comb = 1'h0;
  assign p1_result_i__6_comb = bit_slice_update_w1_1b_1b(p1_result_i__5_comb, p1_result_i__146_comb, p1_result_i__5_comb);
  assign p1_result_i__152_comb = 1'h0;
  assign p1_result_i__15_comb = bit_slice_update_w1_1b_1b(p1_result_i__14_comb, p1_result_i__151_comb, p1_result_i__14_comb);
  assign p1_result_i__157_comb = 1'h0;
  assign p1_result_i__24_comb = bit_slice_update_w1_1b_1b(p1_result_i__23_comb, p1_result_i__156_comb, p1_result_i__23_comb);
  assign p1_result_i__162_comb = 1'h0;
  assign p1_result_i__33_comb = bit_slice_update_w1_1b_1b(p1_result_i__32_comb, p1_result_i__161_comb, p1_result_i__32_comb);
  assign p1_result_i__167_comb = 1'h0;
  assign p1_result_i__42_comb = bit_slice_update_w1_1b_1b(p1_result_i__41_comb, p1_result_i__166_comb, p1_result_i__41_comb);
  assign p1_result_i__172_comb = 1'h0;
  assign p1_result_i__51_comb = bit_slice_update_w1_1b_1b(p1_result_i__50_comb, p1_result_i__171_comb, p1_result_i__50_comb);
  assign p1_result_i__177_comb = 1'h0;
  assign p1_result_i__60_comb = bit_slice_update_w1_1b_1b(p1_result_i__59_comb, p1_result_i__176_comb, p1_result_i__59_comb);
  assign p1_result_i__182_comb = 1'h0;
  assign p1_result_i__69_comb = bit_slice_update_w1_1b_1b(p1_result_i__68_comb, p1_result_i__181_comb, p1_result_i__68_comb);
  assign p1_result_i__187_comb = 1'h0;
  assign p1_result_i__78_comb = bit_slice_update_w1_1b_1b(p1_result_i__77_comb, p1_result_i__186_comb, p1_result_i__77_comb);
  assign p1_result_i__192_comb = 1'h0;
  assign p1_result_i__87_comb = bit_slice_update_w1_1b_1b(p1_result_i__86_comb, p1_result_i__191_comb, p1_result_i__86_comb);
  assign p1_result_i__197_comb = 1'h0;
  assign p1_result_i__96_comb = bit_slice_update_w1_1b_1b(p1_result_i__95_comb, p1_result_i__196_comb, p1_result_i__95_comb);
  assign p1_result_i__202_comb = 1'h0;
  assign p1_result_i__105_comb = bit_slice_update_w1_1b_1b(p1_result_i__104_comb, p1_result_i__201_comb, p1_result_i__104_comb);
  assign p1_result_i__207_comb = 1'h0;
  assign p1_result_i__114_comb = bit_slice_update_w1_1b_1b(p1_result_i__113_comb, p1_result_i__206_comb, p1_result_i__113_comb);
  assign p1_result_i__212_comb = 1'h0;
  assign p1_result_i__123_comb = bit_slice_update_w1_1b_1b(p1_result_i__122_comb, p1_result_i__211_comb, p1_result_i__122_comb);
  assign p1_result_i__217_comb = 1'h0;
  assign p1_result_i__132_comb = bit_slice_update_w1_1b_1b(p1_result_i__131_comb, p1_result_i__216_comb, p1_result_i__131_comb);
  assign p1_result_i__222_comb = 1'h0;
  assign p1_result_i__141_comb = bit_slice_update_w1_1b_1b(p1_result_i__140_comb, p1_result_i__221_comb, p1_result_i__140_comb);
  assign p1_result_i__148_comb = 1'h0;
  assign p1_result_i__7_comb = bit_slice_update_w1_1b_1b(p1_result_i__6_comb, p1_result_i__147_comb, p1_result_i__6_comb);
  assign p1_result_i__153_comb = 1'h0;
  assign p1_result_i__16_comb = bit_slice_update_w1_1b_1b(p1_result_i__15_comb, p1_result_i__152_comb, p1_result_i__15_comb);
  assign p1_result_i__158_comb = 1'h0;
  assign p1_result_i__25_comb = bit_slice_update_w1_1b_1b(p1_result_i__24_comb, p1_result_i__157_comb, p1_result_i__24_comb);
  assign p1_result_i__163_comb = 1'h0;
  assign p1_result_i__34_comb = bit_slice_update_w1_1b_1b(p1_result_i__33_comb, p1_result_i__162_comb, p1_result_i__33_comb);
  assign p1_result_i__168_comb = 1'h0;
  assign p1_result_i__43_comb = bit_slice_update_w1_1b_1b(p1_result_i__42_comb, p1_result_i__167_comb, p1_result_i__42_comb);
  assign p1_result_i__173_comb = 1'h0;
  assign p1_result_i__52_comb = bit_slice_update_w1_1b_1b(p1_result_i__51_comb, p1_result_i__172_comb, p1_result_i__51_comb);
  assign p1_result_i__178_comb = 1'h0;
  assign p1_result_i__61_comb = bit_slice_update_w1_1b_1b(p1_result_i__60_comb, p1_result_i__177_comb, p1_result_i__60_comb);
  assign p1_result_i__183_comb = 1'h0;
  assign p1_result_i__70_comb = bit_slice_update_w1_1b_1b(p1_result_i__69_comb, p1_result_i__182_comb, p1_result_i__69_comb);
  assign p1_result_i__188_comb = 1'h0;
  assign p1_result_i__79_comb = bit_slice_update_w1_1b_1b(p1_result_i__78_comb, p1_result_i__187_comb, p1_result_i__78_comb);
  assign p1_result_i__193_comb = 1'h0;
  assign p1_result_i__88_comb = bit_slice_update_w1_1b_1b(p1_result_i__87_comb, p1_result_i__192_comb, p1_result_i__87_comb);
  assign p1_result_i__198_comb = 1'h0;
  assign p1_result_i__97_comb = bit_slice_update_w1_1b_1b(p1_result_i__96_comb, p1_result_i__197_comb, p1_result_i__96_comb);
  assign p1_result_i__203_comb = 1'h0;
  assign p1_result_i__106_comb = bit_slice_update_w1_1b_1b(p1_result_i__105_comb, p1_result_i__202_comb, p1_result_i__105_comb);
  assign p1_result_i__208_comb = 1'h0;
  assign p1_result_i__115_comb = bit_slice_update_w1_1b_1b(p1_result_i__114_comb, p1_result_i__207_comb, p1_result_i__114_comb);
  assign p1_result_i__213_comb = 1'h0;
  assign p1_result_i__124_comb = bit_slice_update_w1_1b_1b(p1_result_i__123_comb, p1_result_i__212_comb, p1_result_i__123_comb);
  assign p1_result_i__218_comb = 1'h0;
  assign p1_result_i__133_comb = bit_slice_update_w1_1b_1b(p1_result_i__132_comb, p1_result_i__217_comb, p1_result_i__132_comb);
  assign p1_result_i__223_comb = 1'h0;
  assign p1_result_i__142_comb = bit_slice_update_w1_1b_1b(p1_result_i__141_comb, p1_result_i__222_comb, p1_result_i__141_comb);
  assign p1_result_i__8_comb = bit_slice_update_w1_1b_1b(p1_result_i__7_comb, p1_result_i__148_comb, p1_result_i__7_comb);
  assign p1_result_i__17_comb = bit_slice_update_w1_1b_1b(p1_result_i__16_comb, p1_result_i__153_comb, p1_result_i__16_comb);
  assign p1_result_i__26_comb = bit_slice_update_w1_1b_1b(p1_result_i__25_comb, p1_result_i__158_comb, p1_result_i__25_comb);
  assign p1_result_i__35_comb = bit_slice_update_w1_1b_1b(p1_result_i__34_comb, p1_result_i__163_comb, p1_result_i__34_comb);
  assign p1_result_i__44_comb = bit_slice_update_w1_1b_1b(p1_result_i__43_comb, p1_result_i__168_comb, p1_result_i__43_comb);
  assign p1_result_i__53_comb = bit_slice_update_w1_1b_1b(p1_result_i__52_comb, p1_result_i__173_comb, p1_result_i__52_comb);
  assign p1_result_i__62_comb = bit_slice_update_w1_1b_1b(p1_result_i__61_comb, p1_result_i__178_comb, p1_result_i__61_comb);
  assign p1_result_i__71_comb = bit_slice_update_w1_1b_1b(p1_result_i__70_comb, p1_result_i__183_comb, p1_result_i__70_comb);
  assign p1_result_i__80_comb = bit_slice_update_w1_1b_1b(p1_result_i__79_comb, p1_result_i__188_comb, p1_result_i__79_comb);
  assign p1_result_i__89_comb = bit_slice_update_w1_1b_1b(p1_result_i__88_comb, p1_result_i__193_comb, p1_result_i__88_comb);
  assign p1_result_i__98_comb = bit_slice_update_w1_1b_1b(p1_result_i__97_comb, p1_result_i__198_comb, p1_result_i__97_comb);
  assign p1_result_i__107_comb = bit_slice_update_w1_1b_1b(p1_result_i__106_comb, p1_result_i__203_comb, p1_result_i__106_comb);
  assign p1_result_i__116_comb = bit_slice_update_w1_1b_1b(p1_result_i__115_comb, p1_result_i__208_comb, p1_result_i__115_comb);
  assign p1_result_i__125_comb = bit_slice_update_w1_1b_1b(p1_result_i__124_comb, p1_result_i__213_comb, p1_result_i__124_comb);
  assign p1_result_i__134_comb = bit_slice_update_w1_1b_1b(p1_result_i__133_comb, p1_result_i__218_comb, p1_result_i__133_comb);
  assign p1_result_i__143_comb = bit_slice_update_w1_1b_1b(p1_result_i__142_comb, p1_result_i__223_comb, p1_result_i__142_comb);
  assign p1_result__16_comb[0] = p1_result_i__8_comb;
  assign p1_result__16_comb[1] = p1_result_i__17_comb;
  assign p1_result__16_comb[2] = p1_result_i__26_comb;
  assign p1_result__16_comb[3] = p1_result_i__35_comb;
  assign p1_result__16_comb[4] = p1_result_i__44_comb;
  assign p1_result__16_comb[5] = p1_result_i__53_comb;
  assign p1_result__16_comb[6] = p1_result_i__62_comb;
  assign p1_result__16_comb[7] = p1_result_i__71_comb;
  assign p1_result__16_comb[8] = p1_result_i__80_comb;
  assign p1_result__16_comb[9] = p1_result_i__89_comb;
  assign p1_result__16_comb[10] = p1_result_i__98_comb;
  assign p1_result__16_comb[11] = p1_result_i__107_comb;
  assign p1_result__16_comb[12] = p1_result_i__116_comb;
  assign p1_result__16_comb[13] = p1_result_i__125_comb;
  assign p1_result__16_comb[14] = p1_result_i__134_comb;
  assign p1_result__16_comb[15] = p1_result_i__143_comb;

  // Registers for pipe stage 1:
  reg [15:0] p1_result__16;
  always_ff @ (posedge clk) begin
    p1_result__16 <= p1_result__16_comb;
  end
  assign out = {p1_result__16[0], p1_result__16[1], p1_result__16[2], p1_result__16[3], p1_result__16[4], p1_result__16[5], p1_result__16[6], p1_result__16[7], p1_result__16[8], p1_result__16[9], p1_result__16[10], p1_result__16[11], p1_result__16[12], p1_result__16[13], p1_result__16[14], p1_result__16[15]};
endmodule
